library ieee;
use ieee.std_logic_1164.all;

package build_id_pkg is
  constant BUILD_ID : std_logic_vector(31 downto 0) := x"00000000";
end package;
